module get1num_bit(
    input   [7:0]   i_data,
    output  [31:0]  ret
);

endmodule