`ifndef __DEFINE__
`define __DEFINE__


`define DEBUG


`endif